-- TOP LEVEL ENTITY
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY LAB1 IS
	PORT (		
		G_CLOCK_50  : IN  STD_LOGIC;                     -- 50 MHz       (CLOCK)
	
		V_SW        : IN  STD_LOGIC_VECTOR( 7 DOWNTO 0); -- SWITCHES     (A / B)
		V_BT        : IN  STD_LOGIC_VECTOR( 1 DOWNTO 0); -- BUTTONS      (SET / RESET)
		
		G_LEDR		: OUT STD_LOGIC_VECTOR(17 DOWNTO 0); -- RED LEDS     (SWITCHES)
		G_LEDG		: OUT STD_LOGIC_VECTOR( 2 DOWNTO 0); -- GREEN LEDS   (OPT)
		G_HEX7		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (A_1)
		G_HEX6		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (A_0)
		G_HEX5		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (B_1)
		G_HEX4		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (B_0)
		G_HEX3		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (RES_1)
		G_HEX2		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (RES_0)
		G_HEX0		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0)  -- 7SEG DISPLAY (OPT)
		
	);
END LAB1;

ARCHITECTURE BEHAVIORAL OF LAB1 IS
		
	COMPONENT ALU IS  
   PORT (
		A      	: IN   STD_LOGIC_VECTOR(3 DOWNTO 0);
		B      	: IN   STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLK		: IN   STD_LOGIC;
		OPT		: OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		OUTPUT	: OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
   );
	END COMPONENT;
	
	COMPONENT DEC7SEG IS  
   PORT (
		INPUT		: IN   STD_LOGIC_VECTOR(3 DOWNTO 0);
		OUTPUT	: OUT  STD_LOGIC_VECTOR(13 DOWNTO 0)
   );
	END COMPONENT;
	
	COMPONENT FA
	PORT (
		A    : IN  STD_LOGIC;
		B    : IN  STD_LOGIC;
		CIN  : IN  STD_LOGIC;
		S    : OUT STD_LOGIC;
		COUT : OUT STD_LOGIC
	);
	END COMPONENT;
		
	SIGNAL INPUT_A    : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL INPUT_B    : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL INPUT_R    : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL OPT_7SEG   : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL ALU_OPTION : STD_LOGIC_VECTOR( 2 DOWNTO 0);
	SIGNAL ALU_RESULT : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL OUTPUT_A   : STD_LOGIC_VECTOR(13 DOWNTO 0);
	SIGNAL OUTPUT_B   : STD_LOGIC_VECTOR(13 DOWNTO 0);
	SIGNAL OUTPUT_R   : STD_LOGIC_VECTOR(13 DOWNTO 0);
	SIGNAL OUTPUT_OPT : STD_LOGIC_VECTOR(13 DOWNTO 0);
		
	SIGNAL IS_SET     : STD_LOGIC := '0';
	
BEGIN
	
	ALU0: ALU PORT MAP (INPUT_A, INPUT_B, G_CLOCK_50, ALU_OPTION, ALU_RESULT);
	DEC0: DEC7SEG PORT MAP  (INPUT_A,   OUTPUT_A);
	DEC1: DEC7SEG PORT MAP  (INPUT_B,   OUTPUT_B);
	DEC2: DEC7SEG PORT MAP  (INPUT_R,   OUTPUT_R);
	DEC3: DEC7SEG PORT MAP (OPT_7SEG, OUTPUT_OPT);

	PROCESS(INPUT_A, INPUT_B, V_BT, V_SW, OUTPUT_A, OUTPUT_B, OUTPUT_R, OUTPUT_OPT, ALU_RESULT, ALU_OPTION, IS_SET) IS BEGIN
		IF (V_BT(0) = '0') THEN
			IS_SET <= '0';
		ELSIF (V_BT(1) = '0') THEN
			IS_SET <= '1';
		END IF;
		

		IF (IS_SET = '0') THEN
			INPUT_A <= V_SW(7 DOWNTO 4);
			INPUT_B <= V_SW(3 DOWNTO 0);
			INPUT_R <= "0000";
			
			G_LEDR(17 DOWNTO 14) <= INPUT_A;
			G_LEDR(13 DOWNTO 10) <= INPUT_B;
			G_LEDR(3 DOWNTO 0)	<= "0000";
			G_HEX7 <=   OUTPUT_A(13 DOWNTO 7);
			G_HEX6 <=   OUTPUT_A( 6 DOWNTO 0);
			G_HEX5 <=   OUTPUT_B(13 DOWNTO 7);
			G_HEX4 <=   OUTPUT_B( 6 DOWNTO 0);
			G_HEX3 <=   OUTPUT_R(13 DOWNTO 7);
			G_HEX2 <=   OUTPUT_R( 6 DOWNTO 0);
		ELSE
			INPUT_R <= ALU_RESULT;
			
			G_LEDR(3 DOWNTO 0) <= ALU_RESULT;
			G_HEX3 <= OUTPUT_R(13 DOWNTO 7);
			G_HEX2 <= OUTPUT_R( 6 DOWNTO 0);		
		END IF;
		
		OPT_7SEG(2 DOWNTO 0) <= ALU_OPTION;
		G_HEX0 <= OUTPUT_OPT( 6 DOWNTO 0);
		G_LEDG(2 DOWNTO 0) <= ALU_OPTION;
	END PROCESS;
	
END BEHAVIORAL;