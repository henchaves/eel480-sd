-- TOP LEVEL ENTITY
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY LAB2 IS
	PORT (		
		G_CLOCK_50  : IN  STD_LOGIC;                     -- 50 MHz       (CLOCK)
	
		V_SW        : IN  STD_LOGIC_VECTOR(17 DOWNTO 0); -- SWITCHES     (N / OPT)
		V_BT        : IN  STD_LOGIC_VECTOR( 3 DOWNTO 0); -- BUTTONS      (SET A / SET B / -- / RESET)
		
		G_LEDR		: OUT STD_LOGIC_VECTOR(17 DOWNTO 0); -- RED LEDS     (SWITCHES)
		G_LEDG		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- GREEN LEDS   (OPT)
		G_HEX4		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (OPT)
		G_HEX3		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (N_3)
		G_HEX2		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (N_2)
		G_HEX1		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0); -- 7SEG DISPLAY (N_1)
		G_HEX0		: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0)  -- 7SEG DISPLAY (N_0)
		
	);
END LAB2;

ARCHITECTURE BEHAVIORAL OF LAB2 IS
	
	-- 7 SEGMENT DECODER
	COMPONENT DEC7SEG IS  
   PORT (
		INPUT		: IN   STD_LOGIC_VECTOR(3 DOWNTO 0);
		OUTPUT	: OUT  STD_LOGIC_VECTOR(6 DOWNTO 0)
   );
	END COMPONENT;
	
	-- BCD ADDER
	COMPONENT ADDERHANDLER IS
	PORT (
		A    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		S    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
	END COMPONENT;
	
	-- BCD MULTIPLIER
	COMPONENT MULTHANDLER IS
	PORT (
		A    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		P    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
	END COMPONENT;
	
	-- INTERFACE INPUT SIGNALS
	SIGNAL VALUE_A    : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL VALUE_B    : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL VALUE_OPT  : STD_LOGIC := '0';
	
	-- 7 SEGMENT DECODER SIGNALS
	SIGNAL INPUT_0    : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL INPUT_1    : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL INPUT_2    : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL INPUT_3    : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL INPUT_OPT  : STD_LOGIC_VECTOR( 3 DOWNTO 0);
	SIGNAL OUTPUT_0   : STD_LOGIC_VECTOR( 6 DOWNTO 0);
	SIGNAL OUTPUT_1   : STD_LOGIC_VECTOR( 6 DOWNTO 0);
	SIGNAL OUTPUT_2   : STD_LOGIC_VECTOR( 6 DOWNTO 0);
	SIGNAL OUTPUT_3   : STD_LOGIC_VECTOR( 6 DOWNTO 0);
	SIGNAL OUTPUT_OPT : STD_LOGIC_VECTOR( 6 DOWNTO 0);
	
	-- BCD OPERATION SIGNALS
	SIGNAL VALUE_SUM   : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL VALUE_PROD  : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
	
	-- STATE SIGNALS
	SIGNAL SET_A      : STD_LOGIC := '0';
	SIGNAL SET_B      : STD_LOGIC := '0';
	
BEGIN
	
	ADDHAND: ADDERHANDLER PORT MAP (VALUE_A, VALUE_B, VALUE_SUM);
	MULTHAND: MULTHANDLER PORT MAP (VALUE_A, VALUE_B, VALUE_PROD);
	
	DEC0: DEC7SEG PORT MAP   (INPUT_0,   OUTPUT_0);
	DEC1: DEC7SEG PORT MAP   (INPUT_1,   OUTPUT_1);
	DEC2: DEC7SEG PORT MAP   (INPUT_2,   OUTPUT_2);
	DEC3: DEC7SEG PORT MAP   (INPUT_3,   OUTPUT_3);
	DEC4: DEC7SEG PORT MAP (INPUT_OPT, OUTPUT_OPT);

	PROCESS(SET_A, SET_B) IS BEGIN
		-- BUTTON SET_A
		IF ((V_BT(3) = '0') AND (SET_A = '0')) THEN
			SET_A <= '1';
			VALUE_A <= V_SW(17 DOWNTO 2);
		END IF;
		-- BUTTON SET_B
		IF ((V_BT(2) = '0') AND (SET_A = '1') AND (SET_B = '0')) THEN
			SET_B <= '1';
			VALUE_B <= V_SW(17 DOWNTO 2);
		END IF;
		-- BUTTON RESET
		IF (V_BT(0) = '0') THEN
			SET_A <= '0';
			SET_B <= '0';
		END IF;
		
		IF (SET_A = '1') THEN -- IF VALUE_A IS SET
			IF (SET_B = '1') THEN -- IF VALUE_B IS SET
				
				-- BOTH INPUTS ARE SET
				VALUE_OPT <= V_SW(0);
				INPUT_OPT(3 DOWNTO 1) <= "111";
				INPUT_OPT(0) <= VALUE_OPT;
				
				IF (V_SW(0) = '0') THEN -- IF OPT IS SUM
					-- OUTPUTS SUM OF A AND B
					INPUT_0 <= VALUE_SUM( 3 DOWNTO  0);
					INPUT_1 <= VALUE_SUM( 7 DOWNTO  4);
					INPUT_2 <= VALUE_SUM(11 DOWNTO  8);
					INPUT_3 <= VALUE_SUM(15 DOWNTO 12);
					
					G_LEDR <= V_SW;
				ELSE -- IF OPT IS PROD
					-- OUTPUTS PRODUCT OF A AND B
--					INPUT_0(3 DOWNTO 1) <= "111";
--					INPUT_0(0) <= VALUE_OPT;
--					INPUT_1(3 DOWNTO 1) <= "111";
--					INPUT_1(0) <= VALUE_OPT;
--					INPUT_2(3 DOWNTO 1) <= "111";
--					INPUT_2(0) <= VALUE_OPT;
--					INPUT_3(3 DOWNTO 1) <= "111";
--					INPUT_3(0) <= VALUE_OPT;
					INPUT_0 <= VALUE_PROD( 3 DOWNTO  0);
					INPUT_1 <= VALUE_PROD( 7 DOWNTO  4);
					INPUT_2 <= VALUE_PROD(11 DOWNTO  8);
					INPUT_3 <= VALUE_PROD(15 DOWNTO 12);
					
					G_LEDR <= V_SW;
				END IF;
				
			ELSE
				-- ONLY A IS SET
				INPUT_OPT(3 DOWNTO 0) <= "1011";
				INPUT_0 <= V_SW( 5 DOWNTO  2);
				INPUT_1 <= V_SW( 9 DOWNTO  6);
				INPUT_2 <= V_SW(13 DOWNTO 10);
				INPUT_3 <= V_SW(17 DOWNTO 14);
				
				G_LEDR <= V_SW;
			END IF;
		ELSE
			-- NO INPUT IS SET
			INPUT_OPT(3 DOWNTO 0) <= "1010";
			INPUT_0 <= V_SW( 5 DOWNTO  2);
			INPUT_1 <= V_SW( 9 DOWNTO  6);
			INPUT_2 <= V_SW(13 DOWNTO 10);
			INPUT_3 <= V_SW(17 DOWNTO 14);
			
			G_LEDR <= V_SW;
		END IF;
		
		G_LEDG(6) <= SET_A;
		G_LEDG(4) <= SET_B;
		
		G_HEX0 <=   OUTPUT_0( 6 DOWNTO 0);
		G_HEX1 <=   OUTPUT_1( 6 DOWNTO 0);
		G_HEX2 <=   OUTPUT_2( 6 DOWNTO 0);
		G_HEX3 <=   OUTPUT_3( 6 DOWNTO 0);
		G_HEX4 <= OUTPUT_OPT( 6 DOWNTO 0);
		
	END PROCESS;
	
END BEHAVIORAL;