-- 4-BIT BCD ADDER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADDERBCD IS
	PORT (
		A    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		CIN  : IN  STD_LOGIC;
		S    : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		COUT : OUT STD_LOGIC
	);
END ADDERBCD;

ARCHITECTURE BEHAVIORAL OF ADDERBCD IS
	-- 4-BIT BINARY ADDER COMPONENT
	COMPONENT ADDER4BIT
	PORT (
		A    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		CIN  : IN  STD_LOGIC;
		S    : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		COUT : OUT STD_LOGIC
	);
	END COMPONENT;
	
	-- FULL ADDER SIGNALS
	SIGNAL Z      : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL K      : STD_LOGIC;
	SIGNAL OUTC   : STD_LOGIC;
	SIGNAL C      : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL RESULT : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL T      : STD_LOGIC;
BEGIN

	-- FULL ADDER MAPPING
	ADDER4BIT0: ADDER4BIT PORT MAP (A, B, CIN, Z, K);
	ADDER4BIT1: ADDER4BIT PORT MAP (C, Z, '0', RESULT, T);
	
	OUTC <= (K OR (Z(3) AND Z(2)) OR (Z(3) AND Z(1)));
	C(2 DOWNTO 1) <= (OTHERS => OUTC);
	
	S <= RESULT;
	COUT <= OUTC;
	
END BEHAVIORAL;