-- BCD MULTIPLIER HANDLER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ADDERHANDLER IS
	PORT (
		A    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		S    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ADDERHANDLER;

ARCHITECTURE BEHAVIORAL OF ADDERHANDLER IS

	-- 4-BIT BCD ADDER
	COMPONENT ADDERBCD IS
	PORT (
		A    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		CIN  : IN  STD_LOGIC;
		S    : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		COUT : OUT STD_LOGIC
	);
	END COMPONENT;

	-- 4-BIT BCD ADDER SIGNALS
	SIGNAL ADDCOUT0   : STD_LOGIC;
	SIGNAL ADDCOUT1   : STD_LOGIC;
	SIGNAL ADDCOUT2   : STD_LOGIC;
	SIGNAL ADDCOUT3   : STD_LOGIC;
	SIGNAL RESULT     : STD_LOGIC_VECTOR(15 DOWNTO 0);
	
BEGIN
	
	SUM0: ADDERBCD PORT MAP (A( 3 DOWNTO  0), B( 3 DOWNTO  0),      '0', RESULT( 3 DOWNTO  0), ADDCOUT0);
	SUM1: ADDERBCD PORT MAP (A( 7 DOWNTO  4), B( 7 DOWNTO  4), ADDCOUT0, RESULT( 7 DOWNTO  4), ADDCOUT1);
	SUM2: ADDERBCD PORT MAP (A(11 DOWNTO  8), B(11 DOWNTO  8), ADDCOUT1, RESULT(11 DOWNTO  8), ADDCOUT2);
	SUM3: ADDERBCD PORT MAP (A(15 DOWNTO 12), B(15 DOWNTO 12), ADDCOUT2, RESULT(15 DOWNTO 12), ADDCOUT3);
	
	S <= RESULT;
	
		
END BEHAVIORAL;