-- 7SEG BCD DECODER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DEC7SEG IS
	PORT (
		INPUT  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		OUTPUT : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	 );
END ENTITY;
 
ARCHITECTURE BEHAVIORAL OF DEC7SEG IS
BEGIN
	PROCESS(INPUT) IS
	BEGIN
		CASE (INPUT) IS
			WHEN "0000" =>
				OUTPUT <= "10000001000000";
				
			WHEN "0001" =>
				OUTPUT <= "10000001111001";
				
			WHEN "0010" =>
				OUTPUT <= "10000000100100";
				
			WHEN "0011" =>
				OUTPUT <= "10000000110000";
				
			WHEN "0100" =>
				OUTPUT <= "10000000011001";
				
			WHEN "0101" =>
				OUTPUT <= "10000000010010";
				
			WHEN "0110" =>
				OUTPUT <= "10000000000010";
				
			WHEN "0111" =>
				OUTPUT <= "10000001111000";
				
			WHEN "1000" =>
				OUTPUT <= "10000000000000";
				
			WHEN "1001" =>
				OUTPUT <= "10000000010000";
				
			WHEN "1010" =>
				OUTPUT <= "11110011000000";
				
			WHEN "1011" =>
				OUTPUT <= "11110011111001";
				
			WHEN "1100" =>
				OUTPUT <= "11110010100100";
				
			WHEN "1101" =>
				OUTPUT <= "11110010110000";
				
			WHEN "1110" =>
				OUTPUT <= "11110010011001";
				
			WHEN "1111" =>
				OUTPUT <= "11110010010010";
		END CASE;
	END PROCESS;

END ARCHITECTURE;