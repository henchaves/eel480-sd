-- 4x4 MULTIPLIER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MULT IS
	PORT (
		A    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		POUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
	
	SIGNAL C0     : STD_LOGIC := '0';
	SIGNAL C1     : STD_LOGIC := '0';
	SIGNAL C2     : STD_LOGIC := '0';
	SIGNAL C3     : STD_LOGIC := '0';
	SIGNAL TEMP   : STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL PROD   : STD_LOGIC_VECTOR (3 DOWNTO 0);
END MULT;

ARCHITECTURE BEHAVIORAL OF MULT IS
BEGIN

	PROD(0) <= A(0) AND B(0);
	PROD(1) <= (A(1) AND B(0)) XOR (A(0) AND B(1));
	C0 	  <= A(1) AND B(0) AND A(0) AND B(1);
	PROD(2) <= (((A(2) AND B(0)) XOR (A(1) AND B(1))) XOR (A(0) AND B(2))) XOR C0;
	TEMP(0) <= ((A(2) AND B(0)) XOR (A(1) AND B(1)));
	TEMP(1) <= ((A(0) AND B(2)) XOR C0);
	C1 	  <= (A(2) AND B(0) AND A(1) AND B(1));
	C2 	  <= (A(0) AND B(2) AND C0);
	C3 	  <= TEMP(0) AND TEMP(1);
	PROD(3) <= ((((A(3) AND B(0)) XOR (A(2) AND B(1))) XOR (A(1) AND B(2))) XOR (A(0) AND B(3))) XOR C1 XOR C2 XOR C3;
	
	POUT <= PROD;
	
END BEHAVIORAL;