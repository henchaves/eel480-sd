-- 4-BIT BCD MULTIPLIER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MULTBCD IS
	PORT (
		A      : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		B_ALG  : IN  STD_LOGIC_VECTOR( 3 DOWNTO 0);
		FACTOR : IN  INTEGER;
		P      : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END MULTBCD;

ARCHITECTURE BEHAVIORAL OF MULTBCD IS
	
	-- MULTIPLIER SIGNALS
	SIGNAL A_DEC     : INTEGER;
	SIGNAL B_ALG_DEC : INTEGER;
	SIGNAL P_DEC     : INTEGER;
	SIGNAL P0        : INTEGER;
	SIGNAL P1        : INTEGER;
	SIGNAL P2        : INTEGER;
	SIGNAL P3        : INTEGER;
	SIGNAL RESULT    : STD_LOGIC_VECTOR(15 DOWNTO 0);
	
BEGIN
	A_DEC <= TO_INTEGER(UNSIGNED(A(3 DOWNTO 0))) + 10*TO_INTEGER(UNSIGNED(A(7 DOWNTO 4))) + 100*TO_INTEGER(UNSIGNED(A(11 DOWNTO 8))) + 1000*TO_INTEGER(UNSIGNED(A(15 DOWNTO 12)));
	B_ALG_DEC <= TO_INTEGER(UNSIGNED(B_ALG))*FACTOR;
	P_DEC <= A_DEC*B_ALG_DEC;
	
	P0 <= P_DEC MOD 10;
	P1 <= ((P_DEC - P0)/10) MOD 10;
	P2 <= ((P_DEC - P1*10 - P0)/100) MOD 10;
	P3 <= ((P_DEC - P2*100 - P1*10 - P0)/1000) MOD 10;
	
	RESULT( 3 DOWNTO  0) <= STD_LOGIC_VECTOR(TO_UNSIGNED(P0, 4));
	RESULT( 7 DOWNTO  4) <= STD_LOGIC_VECTOR(TO_UNSIGNED(P1, 4));
	RESULT(11 DOWNTO  8) <= STD_LOGIC_VECTOR(TO_UNSIGNED(P2, 4));
	RESULT(15 DOWNTO 12) <= STD_LOGIC_VECTOR(TO_UNSIGNED(P3, 4));
	
	P <= RESULT;
	
		 
END BEHAVIORAL;