-- FULL ADDER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FA IS
	PORT (
		A    : IN  STD_LOGIC;
		B    : IN  STD_LOGIC;
		CIN  : IN  STD_LOGIC;
		S    : OUT STD_LOGIC;
		COUT : OUT STD_LOGIC
	);
END FA;

ARCHITECTURE BEHAVIORAL OF FA IS
BEGIN
	S <= (A XOR B) XOR CIN;
	COUT <= ((A XOR B) AND CIN) OR (A AND B);
END BEHAVIORAL;