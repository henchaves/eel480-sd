-- 4-BIT BINARY ADDER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADDER4BIT IS
	PORT (
		A    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		CIN  : IN  STD_LOGIC;
		S    : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		COUT : OUT STD_LOGIC
	);
END ADDER4BIT;

ARCHITECTURE BEHAVIORAL OF ADDER4BIT IS
	-- FULL ADDER COMPONENT
	COMPONENT FA
	PORT (
		A    : IN  STD_LOGIC;
		B    : IN  STD_LOGIC;
		CIN  : IN  STD_LOGIC;
		S    : OUT STD_LOGIC;
		COUT : OUT STD_LOGIC
	);
	END COMPONENT;
	
	-- FULL ADDER SIGNALS
	SIGNAL FA_C0  : STD_LOGIC := '0';
	SIGNAL FA_C1  : STD_LOGIC := '0';
	SIGNAL FA_C2  : STD_LOGIC := '0';
	SIGNAL FA_C3  : STD_LOGIC := '0';
	SIGNAL FA_OUT : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN

	-- FULL ADDER MAPPING
	FA0: FA PORT MAP (A(0), B(0),    CIN, FA_OUT(0), FA_C0);
	FA1: FA PORT MAP (A(1), B(1),  FA_C0, FA_OUT(1), FA_C1);
	FA2: FA PORT MAP (A(2), B(2),  FA_C1, FA_OUT(2), FA_C2);
	FA3: FA PORT MAP (A(3), B(3),  FA_C2, FA_OUT(3), FA_C3);
	
	S    <= FA_OUT;
	COUT <= FA_C3;
END BEHAVIORAL;