-- 4-BIT BCD MULTIPLIER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.ALL;

ENTITY MULTBCD IS
	PORT (
		A      : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		B_ALG  : IN  STD_LOGIC_VECTOR( 3 DOWNTO 0);
		FACTOR : IN  INTEGER;
		P      : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END MULTBCD;

ARCHITECTURE BEHAVIORAL OF MULTBCD IS
	
	-- MULTIPLIER SIGNALS
	SIGNAL A_DEC     : UNSIGNED;
	SIGNAL B_ALG_DEC : UNSIGNED;
	SIGNAL TEMP      : UNSIGNED;
	SIGNAL P_DEC     : UNSIGNED;
	SIGNAL P0        : UNSIGNED;
	SIGNAL P1        : UNSIGNED;
	SIGNAL P2        : UNSIGNED;
	SIGNAL P3        : UNSIGNED;
	SIGNAL RESULT    : STD_LOGIC_VECTOR(15 DOWNTO 0);
	
BEGIN
	A_DEC <= UNSIGNED(A(3 DOWNTO 0)) + 10*UNSIGNED(A(7 DOWNTO 4)) + 100*UNSIGNED(A(11 DOWNTO 8)) + 1000*UNSIGNED(A(15 DOWNTO 12));
	B_ALG_DEC <= UNSIGNED(B_ALG)*TO_UNSIGNED(FACTOR, B_ALG_DEC'LENGTH);
	P_DEC <= A_DEC*B_ALG_DEC;
	
	P0 <= P_DEC MOD 10;
	P1 <= ((P_DEC - P0)/10) MOD 10;
	P2 <= ((P_DEC - P1*10 - P0)/100) MOD 10;
	P3 <= ((P_DEC - P2*100 - P1*10 - P0)/1000) MOD 10;
	
	RESULT( 3 DOWNTO  0) <= STD_LOGIC_VECTOR(P0)(3 DOWNTO 0);
	RESULT( 7 DOWNTO  4) <= STD_LOGIC_VECTOR(P1)(3 DOWNTO 0);
	RESULT(11 DOWNTO  8) <= STD_LOGIC_VECTOR(P2)(3 DOWNTO 0);
	RESULT(15 DOWNTO 12) <= STD_LOGIC_VECTOR(P3)(3 DOWNTO 0);
	
	P <= RESULT;
	
		 
END BEHAVIORAL;