-- FULL SUBTRACTOR
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FS IS
	PORT (
		A    : IN  STD_LOGIC;
		B    : IN  STD_LOGIC;
		BIN  : IN  STD_LOGIC;
		D    : OUT STD_LOGIC;
		BOUT : OUT STD_LOGIC
	);
END FS;

ARCHITECTURE BEHAVIORAL OF FS IS
BEGIN
	D <= (B XOR BIN) XOR A;
	BOUT <= ((NOT A) AND B) OR ((NOT (A XOR B)) AND BIN);
END BEHAVIORAL;