-- BCD MULTIPLIER HANDLER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MULTHANDLER IS
	PORT (
		A    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		P    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END MULTHANDLER;

ARCHITECTURE BEHAVIORAL OF MULTHANDLER IS
	
	-- 4-BIT BCD MULTIPLIER
	COMPONENT MULTBCD IS
	PORT (
		A      : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		B_ALG  : IN  STD_LOGIC_VECTOR( 3 DOWNTO 0);
		FACTOR : IN  INTEGER;
		P      : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
	END COMPONENT;

	-- BCD ADDER
	COMPONENT ADDERHANDLER IS
	PORT (
		A    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		S    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
	END COMPONENT;
	
	
	-- MULTIPLIER SIGNALS
	SIGNAL MULT0    : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL MULT1    : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL MULT2    : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL MULT3    : STD_LOGIC_VECTOR(15 DOWNTO 0);
	
	-- ADDER SIGNALS
	SIGNAL SUM0     : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL SUM1     : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL SUM2     : STD_LOGIC_VECTOR(15 DOWNTO 0);
	
BEGIN

	MULTBCD0: MULTBCD PORT MAP (A, B( 3 DOWNTO  0), 1, MULT0);
	MULTBCD1: MULTBCD PORT MAP (A, B( 7 DOWNTO  4), 10, MULT1);
	MULTBCD2: MULTBCD PORT MAP (A, B(11 DOWNTO  8), 100, MULT2);
	MULTBCD3: MULTBCD PORT MAP (A, B(15 DOWNTO 12), 1000, MULT3);
	
	ADDHAND0: ADDERHANDLER PORT MAP (MULT0, MULT1, SUM0);
	ADDHAND1: ADDERHANDLER PORT MAP ( SUM0, MULT2, SUM1);
	ADDHAND2: ADDERHANDLER PORT MAP ( SUM1, MULT3, SUM2);
	
	P <= SUM2;
	
		
END BEHAVIORAL;